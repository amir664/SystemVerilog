module Aes_ctr(
    input logic [7:0] nonce[12],
    input logic [7:0] key[32]
);

function return_value name(port_list);
    
endfunction